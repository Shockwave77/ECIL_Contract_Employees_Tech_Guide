----------------------------------------------------------------------------------
-- Company:      ECIL
-- Design Name:  Fundamental Gates
-- Module Name:  Gate_XOR - Behavioral
-- Project Name: 00_Basics
-- Target Devices: Generic FPGA
-- Tool Versions: Any VHDL-2008 compliant tool
-- Description: 
--    Simple 2-input XOR gate.
--    Useful for bit manipulation/parity checks.
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Gate_XOR is
    Port ( 
        a : in  STD_LOGIC;
        b : in  STD_LOGIC;
        y : out STD_LOGIC
    );
end Gate_XOR;

architecture Behavioral of Gate_XOR is
begin
    y <= a xor b;
end Behavioral;
